module state_machine_tb ();

    initial begin
         