module ALU_tb();

    logic[31:0] rs;
    logic[31:0] rt;
    logic[4:0] shift;
    logic[4:0] ALU_ctrl;
    logic[31:0] ALU_out;
    logic[31:0] ALU_lo;
    logic[31:0] ALU_hi;
    logic[2:0] bflag;

    initial begin
        assign rs=10;
        assign rt=7;
        assign ALU_ctrl=0;
        #5 assert(ALU_out==17) else $fatal(1,"Add failed %d",ALU_out);
        assign ALU_ctrl=1;
        #5 assert(ALU_out==3) else $fatal(1,"Sub failed %d",ALU_out);
        assign ALU_ctrl=2;
        assign rs=10;
        assign rt=-7;
        #5 assert(ALU_lo==-70) else $fatal(1,"Mult S lo failed %d",ALU_lo);
        #5 assert(ALU_hi==32'hffffffff) else $fatal(1,"Mult S hi failed %d",ALU_hi);
        assign ALU_ctrl=3;
        assign rs=10;
        assign rt=7;
        #5 assert(ALU_lo==70) else $fatal(1,"Mult US lo failed %d",ALU_lo);
        assert(ALU_hi==32'h00000000) else $fatal(1,"Mult US hi failed %d",ALU_hi);
        assign ALU_ctrl=4;
        assign rs=10;
        assign rt=-2;
        #5 assert(ALU_lo==-5) else $fatal(1,"Div S lo failed %d",ALU_lo);
        assert(ALU_hi==32'hffffffff) else $fatal(1,"Div S hi failed %d",ALU_hi);
        assign ALU_ctrl=5;
        assign rs=21;
        assign rt=4;
        #5 assert(ALU_lo==5) else $fatal(1,"Div US lo failed %d",ALU_lo);
        assert(ALU_hi==0) else $fatal(1,"Div US hi failed %d",ALU_hi);
        assign ALU_ctrl=6;
        assign rs=32'h0A00fff0;
        assign rt=32'h0A0fff00;
        #5 assert(ALU_out==32'h0A00ff00) else $fatal(1,"AND failed %d",ALU_out);
        assign ALU_ctrl=7;
        assign rs=32'h0A00fff0;
        assign rt=32'h0A0fff00;
        #5 assert(ALU_out==32'h0A0ffff0) else $fatal(1,"OR failed %d",ALU_out);
        assign ALU_ctrl=8;
        assign rs=32'h0A00fff0;
        assign rt=32'h0A0fff00;
        #5 assert(ALU_out==32'h000f00f0) else $fatal(1,"XOR failed %d",ALU_out);
        assign ALU_ctrl=9;
        assign rs=32'h0A00fff0;
        assign rt=32'h00000A08;
        assign shift=4;
        #5 assert(ALU_out==32'hA00fff00) else $fatal(1,"SLL failed %d",ALU_out);
        assign ALU_ctrl=10;
        #5 assert(ALU_out==32'h00fff000) else $fatal(1,"SLV failed %d",ALU_out);
        assign ALU_ctrl=11;
        assign rs=32'h0A00fff0;
        assign rt=32'h00000A08;
        assign shift=4;
        #5 assert(ALU_out==32'h00A00fff) else $fatal(1,"SRL failed %d",ALU_out);
        assign ALU_ctrl=12;
        #5 assert(ALU_out==32'h000A00ff) else $fatal(1,"SRLV failed %d",ALU_out);
        assign ALU_ctrl=13;
        assign rs=32'hfA00fff0;
        assign rt=32'h00000A08;
        assign shift=4;
        #5 assert(ALU_out==32'hffA00fff) else $fatal(1,"SRA failed %d",ALU_out);
        assign ALU_ctrl=14;
        assign rs=32'hAA00fff0;
        #5 assert(ALU_out==32'hffAA00ff) else $fatal(1,"SRAV failed %d",ALU_out);
        assign ALU_ctrl=15;
        assign rs=12;
        assign rt=12;
        #5 assert(ALU_out==1) else $fatal(1,"equals failed %d",ALU_out);
        #5 assert(bflag==0) else $fatal(1,"equals failed %d",bflag);
        assign rt=13;
        #5 assert(ALU_out==0) else $fatal(1,"equals failed %d",ALU_out);
        assign ALU_ctrl=16;
        assign rs=12;
        #5 assert(ALU_out==1) else $fatal(1,"gez failed %d",ALU_out);
        #5 assert(bflag==1) else $fatal(1,"gez failed %d",bflag);
        assign rs=-1;
        #5 assert(ALU_out==0) else $fatal(1,"gez failed %d",ALU_out);
        assign ALU_ctrl=17;
        assign rs=12;
        #5 assert(ALU_out==1) else $fatal(1,"gz failed %d",ALU_out);
        #5 assert(bflag==2) else $fatal(1,"gz failed %d",bflag);
        assign rs=0;
        #5 assert(ALU_out==0) else $fatal(1,"gz failed %d",ALU_out);
        assign ALU_ctrl=18;
        assign rs=-12;
        #5 assert(ALU_out==1) else $fatal(1,"lez failed %d",ALU_out);
        #5 assert(bflag==3) else $fatal(1,"lez failed %d",bflag);
        assign rs=1;
        #5 assert(ALU_out==0) else $fatal(1,"lez failed %d",ALU_out);
        assign ALU_ctrl=19;
        assign rs=-12;
        #5 assert(ALU_out==1) else $fatal(1,"lz failed %d",ALU_out);
        #5 assert(bflag==4) else $fatal(1,"lz failed %d",bflag);
        assign rs=0;
        #5 assert(ALU_out==0) else $fatal(1,"lz failed %d",ALU_out);
        assign ALU_ctrl=20;
        assign rs=12;
        assign rt=10;
        #5 assert(ALU_out==1) else $fatal(1,"ne failed %d",ALU_out);
        #5 assert(bflag==5) else $fatal(1,"ne failed %d",bflag);
        assign rs=10;
        #5 assert(ALU_out==0) else $fatal(1,"ne failed %d",ALU_out);


    end

    ALU dut(rs, rt, shift, ALU_ctrl, ALU_out, ALU_lo, ALU_hi, bflag);

endmodule