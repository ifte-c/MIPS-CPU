module control(
    input logic[5:0] op,
    output logic
);