module decoder(
    logic[31:0] instr,
    
);